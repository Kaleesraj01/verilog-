// dataflow 
module basic_gates(input a,b,output and_out,or_out);
assign and_out= a&b;
assign or_out= a|b;
endmodule
