module and_gate(input a,b,output c );
and (c,a,b);
endmodule

